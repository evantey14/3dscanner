`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    17:42:00 11/27/2016 
// Design Name: 
// Module Name:    write_to_zbt 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module manual_write_to_zbt(
	input clk,
	input [18:0] size,
	output reg [18+2:0] addr,
	output reg [35:0] value
    );
	
	 always @(posedge clk) begin
		if (addr[20:2] > size) addr <= 0;
		else addr <= addr+1;
	 end
	 
	 always @(addr)
		case (addr)
	7'd0: value = {6'b0,-10'd100,-10'd100,-10'd100};
	7'd1: value = {6'b0,-10'd100,-10'd100,-10'd50};
	7'd2: value = {6'b0,-10'd100,-10'd100,10'd0};
	7'd3: value = {6'b0,-10'd100,-10'd100,10'd50};
	7'd4: value = {6'b0,-10'd100,-10'd100,10'd100};
	7'd5: value = {6'b0,-10'd100,-10'd50,-10'd100};
	7'd6: value = {6'b0,-10'd100,-10'd50,-10'd50};
	7'd7: value = {6'b0,-10'd100,-10'd50,10'd0};
	7'd8: value = {6'b0,-10'd100,-10'd50,10'd50};
	7'd9: value = {6'b0,-10'd100,-10'd50,10'd100};
	7'd10: value = {6'b0,-10'd100,10'd0,-10'd100};
	7'd11: value = {6'b0,-10'd100,10'd0,-10'd50};
	7'd12: value = {6'b0,-10'd100,10'd0,10'd0};
	7'd13: value = {6'b0,-10'd100,10'd0,10'd50};
	7'd14: value = {6'b0,-10'd100,10'd0,10'd100};
	7'd15: value = {6'b0,-10'd100,10'd50,-10'd100};
	7'd16: value = {6'b0,-10'd100,10'd50,-10'd50};
	7'd17: value = {6'b0,-10'd100,10'd50,10'd0};
	7'd18: value = {6'b0,-10'd100,10'd50,10'd50};
	7'd19: value = {6'b0,-10'd100,10'd50,10'd100};
	7'd20: value = {6'b0,-10'd100,10'd100,-10'd100};
	7'd21: value = {6'b0,-10'd100,10'd100,-10'd50};
	7'd22: value = {6'b0,-10'd100,10'd100,10'd0};
	7'd23: value = {6'b0,-10'd100,10'd100,10'd50};
	7'd24: value = {6'b0,-10'd100,10'd100,10'd100};
	7'd25: value = {6'b0,-10'd50,-10'd100,-10'd100};
	7'd26: value = {6'b0,-10'd50,-10'd100,-10'd50};
	7'd27: value = {6'b0,-10'd50,-10'd100,10'd0};
	7'd28: value = {6'b0,-10'd50,-10'd100,10'd50};
	7'd29: value = {6'b0,-10'd50,-10'd100,10'd100};
	7'd30: value = {6'b0,-10'd50,-10'd50,-10'd100};
	7'd31: value = {6'b0,-10'd50,-10'd50,-10'd50};
	7'd32: value = {6'b0,-10'd50,-10'd50,10'd0};
	7'd33: value = {6'b0,-10'd50,-10'd50,10'd50};
	7'd34: value = {6'b0,-10'd50,-10'd50,10'd100};
	7'd35: value = {6'b0,-10'd50,10'd0,-10'd100};
	7'd36: value = {6'b0,-10'd50,10'd0,-10'd50};
	7'd37: value = {6'b0,-10'd50,10'd0,10'd0};
	7'd38: value = {6'b0,-10'd50,10'd0,10'd50};
	7'd39: value = {6'b0,-10'd50,10'd0,10'd100};
	7'd40: value = {6'b0,-10'd50,10'd50,-10'd100};
	7'd41: value = {6'b0,-10'd50,10'd50,-10'd50};
	7'd42: value = {6'b0,-10'd50,10'd50,10'd0};
	7'd43: value = {6'b0,-10'd50,10'd50,10'd50};
	7'd44: value = {6'b0,-10'd50,10'd50,10'd100};
	7'd45: value = {6'b0,-10'd50,10'd100,-10'd100};
	7'd46: value = {6'b0,-10'd50,10'd100,-10'd50};
	7'd47: value = {6'b0,-10'd50,10'd100,10'd0};
	7'd48: value = {6'b0,-10'd50,10'd100,10'd50};
	7'd49: value = {6'b0,-10'd50,10'd100,10'd100};
	7'd50: value = {6'b0,10'd0,-10'd100,-10'd100};
	7'd51: value = {6'b0,10'd0,-10'd100,-10'd50};
	7'd52: value = {6'b0,10'd0,-10'd100,10'd0};
	7'd53: value = {6'b0,10'd0,-10'd100,10'd50};
	7'd54: value = {6'b0,10'd0,-10'd100,10'd100};
	7'd55: value = {6'b0,10'd0,-10'd50,-10'd100};
	7'd56: value = {6'b0,10'd0,-10'd50,-10'd50};
	7'd57: value = {6'b0,10'd0,-10'd50,10'd0};
	7'd58: value = {6'b0,10'd0,-10'd50,10'd50};
	7'd59: value = {6'b0,10'd0,-10'd50,10'd100};
	7'd60: value = {6'b0,10'd0,10'd0,-10'd100};
	7'd61: value = {6'b0,10'd0,10'd0,-10'd50};
	7'd62: value = {6'b0,10'd0,10'd0,10'd0};
	7'd63: value = {6'b0,10'd0,10'd0,10'd50};
	7'd64: value = {6'b0,10'd0,10'd0,10'd100};
	7'd65: value = {6'b0,10'd0,10'd50,-10'd100};
	7'd66: value = {6'b0,10'd0,10'd50,-10'd50};
	7'd67: value = {6'b0,10'd0,10'd50,10'd0};
	7'd68: value = {6'b0,10'd0,10'd50,10'd50};
	7'd69: value = {6'b0,10'd0,10'd50,10'd100};
	7'd70: value = {6'b0,10'd0,10'd100,-10'd100};
	7'd71: value = {6'b0,10'd0,10'd100,-10'd50};
	7'd72: value = {6'b0,10'd0,10'd100,10'd0};
	7'd73: value = {6'b0,10'd0,10'd100,10'd50};
	7'd74: value = {6'b0,10'd0,10'd100,10'd100};
	7'd75: value = {6'b0,10'd50,-10'd100,-10'd100};
	7'd76: value = {6'b0,10'd50,-10'd100,-10'd50};
	7'd77: value = {6'b0,10'd50,-10'd100,10'd0};
	7'd78: value = {6'b0,10'd50,-10'd100,10'd50};
	7'd79: value = {6'b0,10'd50,-10'd100,10'd100};
	7'd80: value = {6'b0,10'd50,-10'd50,-10'd100};
	7'd81: value = {6'b0,10'd50,-10'd50,-10'd50};
	7'd82: value = {6'b0,10'd50,-10'd50,10'd0};
	7'd83: value = {6'b0,10'd50,-10'd50,10'd50};
	7'd84: value = {6'b0,10'd50,-10'd50,10'd100};
	7'd85: value = {6'b0,10'd50,10'd0,-10'd100};
	7'd86: value = {6'b0,10'd50,10'd0,-10'd50};
	7'd87: value = {6'b0,10'd50,10'd0,10'd0};
	7'd88: value = {6'b0,10'd50,10'd0,10'd50};
	7'd89: value = {6'b0,10'd50,10'd0,10'd100};
	7'd90: value = {6'b0,10'd50,10'd50,-10'd100};
	7'd91: value = {6'b0,10'd50,10'd50,-10'd50};
	7'd92: value = {6'b0,10'd50,10'd50,10'd0};
	7'd93: value = {6'b0,10'd50,10'd50,10'd50};
	7'd94: value = {6'b0,10'd50,10'd50,10'd100};
	7'd95: value = {6'b0,10'd50,10'd100,-10'd100};
	7'd96: value = {6'b0,10'd50,10'd100,-10'd50};
	7'd97: value = {6'b0,10'd50,10'd100,10'd0};
	7'd98: value = {6'b0,10'd50,10'd100,10'd50};
	7'd99: value = {6'b0,10'd50,10'd100,10'd100};
	7'd100: value = {6'b0,10'd100,-10'd100,-10'd100};
	7'd101: value = {6'b0,10'd100,-10'd100,-10'd50};
	7'd102: value = {6'b0,10'd100,-10'd100,10'd0};
	7'd103: value = {6'b0,10'd100,-10'd100,10'd50};
	7'd104: value = {6'b0,10'd100,-10'd100,10'd100};
	7'd105: value = {6'b0,10'd100,-10'd50,-10'd100};
	7'd106: value = {6'b0,10'd100,-10'd50,-10'd50};
	7'd107: value = {6'b0,10'd100,-10'd50,10'd0};
	7'd108: value = {6'b0,10'd100,-10'd50,10'd50};
	7'd109: value = {6'b0,10'd100,-10'd50,10'd100};
	7'd110: value = {6'b0,10'd100,10'd0,-10'd100};
	7'd111: value = {6'b0,10'd100,10'd0,-10'd50};
	7'd112: value = {6'b0,10'd100,10'd0,10'd0};
	7'd113: value = {6'b0,10'd100,10'd0,10'd50};
	7'd114: value = {6'b0,10'd100,10'd0,10'd100};
	7'd115: value = {6'b0,10'd100,10'd50,-10'd100};
	7'd116: value = {6'b0,10'd100,10'd50,-10'd50};
	7'd117: value = {6'b0,10'd100,10'd50,10'd0};
	7'd118: value = {6'b0,10'd100,10'd50,10'd50};
	7'd119: value = {6'b0,10'd100,10'd50,10'd100};
	7'd120: value = {6'b0,10'd100,10'd100,-10'd100};
	7'd121: value = {6'b0,10'd100,10'd100,-10'd50};
	7'd122: value = {6'b0,10'd100,10'd100,10'd0};
	7'd123: value = {6'b0,10'd100,10'd100,10'd50};
	7'd124: value = {6'b0,10'd100,10'd100,10'd100};
	7'd125: value = {6'b0,10'd200,10'd100,10'd100};
	7'd126: value = {6'b0,10'd200,-10'd100,10'd100};
	7'd127: value = {6'b0,10'd200,10'd100,-10'd100};
			default: value = 0;
		endcase
endmodule
