`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    17:42:00 11/27/2016 
// Design Name: 
// Module Name:    write_to_zbt 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module write_to_zbt(
	input wire [8:0] index,
	output reg [35:0] value
    );
	 always @(index)
		case (index)
			9'd0: value = {6'b0,-10'd0,-10'd58,-10'd341};
9'd1: value = {6'b0,-10'd0,-10'd93,-10'd306};
9'd2: value = {6'b0,-10'd0,-10'd129,-10'd270};
9'd3: value = {6'b0,-10'd0,-10'd164,-10'd235};
9'd4: value = {6'b0,-10'd0,-10'd200,-10'd199};
9'd5: value = {6'b0,-10'd0,-10'd235,-10'd164};
9'd6: value = {6'b0,-10'd0,-10'd270,-10'd129};
9'd7: value = {6'b0,-10'd0,-10'd306,-10'd93};
9'd8: value = {6'b0,-10'd35,-10'd33,-10'd316};
9'd9: value = {6'b0,-10'd35,-10'd68,-10'd281};
9'd10: value = {6'b0,-10'd35,-10'd104,-10'd245};
9'd11: value = {6'b0,-10'd35,-10'd139,-10'd210};
9'd12: value = {6'b0,-10'd35,-10'd175,-10'd174};
9'd13: value = {6'b0,-10'd35,-10'd210,-10'd139};
9'd14: value = {6'b0,-10'd35,-10'd245,-10'd104};
9'd15: value = {6'b0,-10'd35,-10'd281,-10'd68};
9'd16: value = {6'b0,-10'd70,-10'd8,-10'd291};
9'd17: value = {6'b0,-10'd70,-10'd43,-10'd256};
9'd18: value = {6'b0,-10'd70,-10'd79,-10'd220};
9'd19: value = {6'b0,-10'd70,-10'd114,-10'd185};
9'd20: value = {6'b0,-10'd70,-10'd150,-10'd149};
9'd21: value = {6'b0,-10'd70,-10'd185,-10'd114};
9'd22: value = {6'b0,-10'd70,-10'd220,-10'd79};
9'd23: value = {6'b0,-10'd70,-10'd256,-10'd43};
9'd24: value = {6'b0,-10'd106,10'd16,-10'd266};
9'd25: value = {6'b0,-10'd106,-10'd18,-10'd231};
9'd26: value = {6'b0,-10'd106,-10'd54,-10'd195};
9'd27: value = {6'b0,-10'd106,-10'd89,-10'd160};
9'd28: value = {6'b0,-10'd106,-10'd125,-10'd124};
9'd29: value = {6'b0,-10'd106,-10'd160,-10'd89};
9'd30: value = {6'b0,-10'd106,-10'd195,-10'd54};
9'd31: value = {6'b0,-10'd106,-10'd231,-10'd18};
9'd32: value = {6'b0,-10'd141,10'd41,-10'd241};
9'd33: value = {6'b0,-10'd141,10'd6,-10'd206};
9'd34: value = {6'b0,-10'd141,-10'd29,-10'd170};
9'd35: value = {6'b0,-10'd141,-10'd64,-10'd135};
9'd36: value = {6'b0,-10'd141,-10'd99,-10'd99};
9'd37: value = {6'b0,-10'd141,-10'd135,-10'd64};
9'd38: value = {6'b0,-10'd141,-10'd170,-10'd29};
9'd39: value = {6'b0,-10'd141,-10'd206,10'd6};
9'd40: value = {6'b0,-10'd176,10'd66,-10'd216};
9'd41: value = {6'b0,-10'd176,10'd31,-10'd181};
9'd42: value = {6'b0,-10'd176,-10'd4,-10'd145};
9'd43: value = {6'b0,-10'd176,-10'd39,-10'd110};
9'd44: value = {6'b0,-10'd176,-10'd74,-10'd74};
9'd45: value = {6'b0,-10'd176,-10'd110,-10'd39};
9'd46: value = {6'b0,-10'd176,-10'd145,-10'd4};
9'd47: value = {6'b0,-10'd176,-10'd181,10'd31};
9'd48: value = {6'b0,-10'd212,10'd91,-10'd191};
9'd49: value = {6'b0,-10'd212,10'd56,-10'd156};
9'd50: value = {6'b0,-10'd212,10'd20,-10'd120};
9'd51: value = {6'b0,-10'd212,-10'd14,-10'd85};
9'd52: value = {6'b0,-10'd212,-10'd49,-10'd49};
9'd53: value = {6'b0,-10'd212,-10'd85,-10'd14};
9'd54: value = {6'b0,-10'd212,-10'd120,10'd20};
9'd55: value = {6'b0,-10'd212,-10'd156,10'd56};
9'd56: value = {6'b0,-10'd247,10'd116,-10'd166};
9'd57: value = {6'b0,-10'd247,10'd81,-10'd131};
9'd58: value = {6'b0,-10'd247,10'd45,-10'd95};
9'd59: value = {6'b0,-10'd247,10'd10,-10'd60};
9'd60: value = {6'b0,-10'd247,-10'd24,-10'd24};
9'd61: value = {6'b0,-10'd247,-10'd60,10'd10};
9'd62: value = {6'b0,-10'd247,-10'd95,10'd45};
9'd63: value = {6'b0,-10'd247,-10'd131,10'd81};
9'd64: value = {6'b0,10'd35,-10'd33,-10'd316};
9'd65: value = {6'b0,10'd35,-10'd68,-10'd281};
9'd66: value = {6'b0,10'd35,-10'd104,-10'd245};
9'd67: value = {6'b0,10'd35,-10'd139,-10'd210};
9'd68: value = {6'b0,10'd35,-10'd175,-10'd174};
9'd69: value = {6'b0,10'd35,-10'd210,-10'd139};
9'd70: value = {6'b0,10'd35,-10'd245,-10'd104};
9'd71: value = {6'b0,10'd35,-10'd281,-10'd68};
9'd72: value = {6'b0,-10'd0,-10'd8,-10'd291};
9'd73: value = {6'b0,-10'd0,-10'd43,-10'd256};
9'd74: value = {6'b0,-10'd0,-10'd79,-10'd220};
9'd75: value = {6'b0,-10'd0,-10'd114,-10'd185};
9'd76: value = {6'b0,-10'd0,-10'd150,-10'd149};
9'd77: value = {6'b0,-10'd0,-10'd185,-10'd114};
9'd78: value = {6'b0,-10'd0,-10'd220,-10'd79};
9'd79: value = {6'b0,-10'd0,-10'd256,-10'd43};
9'd80: value = {6'b0,-10'd35,10'd16,-10'd266};
9'd81: value = {6'b0,-10'd35,-10'd18,-10'd231};
9'd82: value = {6'b0,-10'd35,-10'd54,-10'd195};
9'd83: value = {6'b0,-10'd35,-10'd89,-10'd160};
9'd84: value = {6'b0,-10'd35,-10'd125,-10'd124};
9'd85: value = {6'b0,-10'd35,-10'd160,-10'd89};
9'd86: value = {6'b0,-10'd35,-10'd195,-10'd54};
9'd87: value = {6'b0,-10'd35,-10'd231,-10'd18};
9'd88: value = {6'b0,-10'd70,10'd41,-10'd241};
9'd89: value = {6'b0,-10'd70,10'd6,-10'd206};
9'd90: value = {6'b0,-10'd70,-10'd29,-10'd170};
9'd91: value = {6'b0,-10'd70,-10'd64,-10'd135};
9'd92: value = {6'b0,-10'd70,-10'd100,-10'd99};
9'd93: value = {6'b0,-10'd70,-10'd135,-10'd64};
9'd94: value = {6'b0,-10'd70,-10'd170,-10'd29};
9'd95: value = {6'b0,-10'd70,-10'd206,10'd6};
9'd96: value = {6'b0,-10'd106,10'd66,-10'd216};
9'd97: value = {6'b0,-10'd106,10'd31,-10'd181};
9'd98: value = {6'b0,-10'd106,-10'd4,-10'd145};
9'd99: value = {6'b0,-10'd106,-10'd39,-10'd110};
9'd100: value = {6'b0,-10'd106,-10'd74,-10'd74};
9'd101: value = {6'b0,-10'd106,-10'd110,-10'd39};
9'd102: value = {6'b0,-10'd106,-10'd145,-10'd4};
9'd103: value = {6'b0,-10'd106,-10'd181,10'd31};
9'd104: value = {6'b0,-10'd141,10'd91,-10'd191};
9'd105: value = {6'b0,-10'd141,10'd56,-10'd156};
9'd106: value = {6'b0,-10'd141,10'd20,-10'd120};
9'd107: value = {6'b0,-10'd141,-10'd14,-10'd85};
9'd108: value = {6'b0,-10'd141,-10'd49,-10'd49};
9'd109: value = {6'b0,-10'd141,-10'd85,-10'd14};
9'd110: value = {6'b0,-10'd141,-10'd120,10'd20};
9'd111: value = {6'b0,-10'd141,-10'd156,10'd56};
9'd112: value = {6'b0,-10'd176,10'd116,-10'd166};
9'd113: value = {6'b0,-10'd176,10'd81,-10'd131};
9'd114: value = {6'b0,-10'd176,10'd45,-10'd95};
9'd115: value = {6'b0,-10'd176,10'd10,-10'd60};
9'd116: value = {6'b0,-10'd176,-10'd24,-10'd24};
9'd117: value = {6'b0,-10'd176,-10'd60,10'd10};
9'd118: value = {6'b0,-10'd176,-10'd95,10'd45};
9'd119: value = {6'b0,-10'd176,-10'd131,10'd81};
9'd120: value = {6'b0,-10'd212,10'd141,-10'd141};
9'd121: value = {6'b0,-10'd212,10'd106,-10'd106};
9'd122: value = {6'b0,-10'd212,10'd70,-10'd70};
9'd123: value = {6'b0,-10'd212,10'd35,-10'd35};
9'd124: value = {6'b0,-10'd212,10'd0,10'd0};
9'd125: value = {6'b0,-10'd212,-10'd35,10'd35};
9'd126: value = {6'b0,-10'd212,-10'd70,10'd70};
9'd127: value = {6'b0,-10'd212,-10'd106,10'd106};
9'd128: value = {6'b0,10'd70,-10'd8,-10'd291};
9'd129: value = {6'b0,10'd70,-10'd43,-10'd256};
9'd130: value = {6'b0,10'd70,-10'd79,-10'd220};
9'd131: value = {6'b0,10'd70,-10'd114,-10'd185};
9'd132: value = {6'b0,10'd70,-10'd150,-10'd149};
9'd133: value = {6'b0,10'd70,-10'd185,-10'd114};
9'd134: value = {6'b0,10'd70,-10'd220,-10'd79};
9'd135: value = {6'b0,10'd70,-10'd256,-10'd43};
9'd136: value = {6'b0,10'd35,10'd16,-10'd266};
9'd137: value = {6'b0,10'd35,-10'd18,-10'd231};
9'd138: value = {6'b0,10'd35,-10'd54,-10'd195};
9'd139: value = {6'b0,10'd35,-10'd89,-10'd160};
9'd140: value = {6'b0,10'd35,-10'd125,-10'd124};
9'd141: value = {6'b0,10'd35,-10'd160,-10'd89};
9'd142: value = {6'b0,10'd35,-10'd195,-10'd54};
9'd143: value = {6'b0,10'd35,-10'd231,-10'd18};
9'd144: value = {6'b0,-10'd0,10'd41,-10'd241};
9'd145: value = {6'b0,-10'd0,10'd6,-10'd206};
9'd146: value = {6'b0,-10'd0,-10'd29,-10'd170};
9'd147: value = {6'b0,-10'd0,-10'd64,-10'd135};
9'd148: value = {6'b0,-10'd0,-10'd100,-10'd99};
9'd149: value = {6'b0,-10'd0,-10'd135,-10'd64};
9'd150: value = {6'b0,-10'd0,-10'd170,-10'd29};
9'd151: value = {6'b0,-10'd0,-10'd206,10'd6};
9'd152: value = {6'b0,-10'd35,10'd66,-10'd216};
9'd153: value = {6'b0,-10'd35,10'd31,-10'd181};
9'd154: value = {6'b0,-10'd35,-10'd4,-10'd145};
9'd155: value = {6'b0,-10'd35,-10'd39,-10'd110};
9'd156: value = {6'b0,-10'd35,-10'd75,-10'd74};
9'd157: value = {6'b0,-10'd35,-10'd110,-10'd39};
9'd158: value = {6'b0,-10'd35,-10'd145,-10'd4};
9'd159: value = {6'b0,-10'd35,-10'd181,10'd31};
9'd160: value = {6'b0,-10'd70,10'd91,-10'd191};
9'd161: value = {6'b0,-10'd70,10'd56,-10'd156};
9'd162: value = {6'b0,-10'd70,10'd20,-10'd120};
9'd163: value = {6'b0,-10'd70,-10'd14,-10'd85};
9'd164: value = {6'b0,-10'd70,-10'd49,-10'd49};
9'd165: value = {6'b0,-10'd70,-10'd85,-10'd14};
9'd166: value = {6'b0,-10'd70,-10'd120,10'd20};
9'd167: value = {6'b0,-10'd70,-10'd156,10'd56};
9'd168: value = {6'b0,-10'd106,10'd116,-10'd166};
9'd169: value = {6'b0,-10'd106,10'd81,-10'd131};
9'd170: value = {6'b0,-10'd106,10'd45,-10'd95};
9'd171: value = {6'b0,-10'd106,10'd10,-10'd60};
9'd172: value = {6'b0,-10'd106,-10'd24,-10'd24};
9'd173: value = {6'b0,-10'd106,-10'd60,10'd10};
9'd174: value = {6'b0,-10'd106,-10'd95,10'd45};
9'd175: value = {6'b0,-10'd106,-10'd131,10'd81};
9'd176: value = {6'b0,-10'd141,10'd141,-10'd141};
9'd177: value = {6'b0,-10'd141,10'd106,-10'd106};
9'd178: value = {6'b0,-10'd141,10'd70,-10'd70};
9'd179: value = {6'b0,-10'd141,10'd35,-10'd35};
9'd180: value = {6'b0,-10'd141,10'd0,10'd0};
9'd181: value = {6'b0,-10'd141,-10'd35,10'd35};
9'd182: value = {6'b0,-10'd141,-10'd70,10'd70};
9'd183: value = {6'b0,-10'd141,-10'd106,10'd106};
9'd184: value = {6'b0,-10'd176,10'd166,-10'd116};
9'd185: value = {6'b0,-10'd176,10'd131,-10'd81};
9'd186: value = {6'b0,-10'd176,10'd95,-10'd45};
9'd187: value = {6'b0,-10'd176,10'd60,-10'd10};
9'd188: value = {6'b0,-10'd176,10'd25,10'd25};
9'd189: value = {6'b0,-10'd176,-10'd10,10'd60};
9'd190: value = {6'b0,-10'd176,-10'd45,10'd95};
9'd191: value = {6'b0,-10'd176,-10'd81,10'd131};
9'd192: value = {6'b0,10'd106,10'd16,-10'd266};
9'd193: value = {6'b0,10'd106,-10'd18,-10'd231};
9'd194: value = {6'b0,10'd106,-10'd54,-10'd195};
9'd195: value = {6'b0,10'd106,-10'd89,-10'd160};
9'd196: value = {6'b0,10'd106,-10'd125,-10'd124};
9'd197: value = {6'b0,10'd106,-10'd160,-10'd89};
9'd198: value = {6'b0,10'd106,-10'd195,-10'd54};
9'd199: value = {6'b0,10'd106,-10'd231,-10'd18};
9'd200: value = {6'b0,10'd70,10'd41,-10'd241};
9'd201: value = {6'b0,10'd70,10'd6,-10'd206};
9'd202: value = {6'b0,10'd70,-10'd29,-10'd170};
9'd203: value = {6'b0,10'd70,-10'd64,-10'd135};
9'd204: value = {6'b0,10'd70,-10'd100,-10'd99};
9'd205: value = {6'b0,10'd70,-10'd135,-10'd64};
9'd206: value = {6'b0,10'd70,-10'd170,-10'd29};
9'd207: value = {6'b0,10'd70,-10'd206,10'd6};
9'd208: value = {6'b0,10'd35,10'd66,-10'd216};
9'd209: value = {6'b0,10'd35,10'd31,-10'd181};
9'd210: value = {6'b0,10'd35,-10'd4,-10'd145};
9'd211: value = {6'b0,10'd35,-10'd39,-10'd110};
9'd212: value = {6'b0,10'd35,-10'd75,-10'd74};
9'd213: value = {6'b0,10'd35,-10'd110,-10'd39};
9'd214: value = {6'b0,10'd35,-10'd145,-10'd4};
9'd215: value = {6'b0,10'd35,-10'd181,10'd31};
9'd216: value = {6'b0,-10'd0,10'd91,-10'd191};
9'd217: value = {6'b0,-10'd0,10'd56,-10'd156};
9'd218: value = {6'b0,-10'd0,10'd20,-10'd120};
9'd219: value = {6'b0,-10'd0,-10'd14,-10'd85};
9'd220: value = {6'b0,-10'd0,-10'd50,-10'd49};
9'd221: value = {6'b0,-10'd0,-10'd85,-10'd14};
9'd222: value = {6'b0,-10'd0,-10'd120,10'd20};
9'd223: value = {6'b0,-10'd0,-10'd156,10'd56};
9'd224: value = {6'b0,-10'd35,10'd116,-10'd166};
9'd225: value = {6'b0,-10'd35,10'd81,-10'd131};
9'd226: value = {6'b0,-10'd35,10'd45,-10'd95};
9'd227: value = {6'b0,-10'd35,10'd10,-10'd60};
9'd228: value = {6'b0,-10'd35,-10'd24,-10'd24};
9'd229: value = {6'b0,-10'd35,-10'd60,10'd10};
9'd230: value = {6'b0,-10'd35,-10'd95,10'd45};
9'd231: value = {6'b0,-10'd35,-10'd131,10'd81};
9'd232: value = {6'b0,-10'd70,10'd141,-10'd141};
9'd233: value = {6'b0,-10'd70,10'd106,-10'd106};
9'd234: value = {6'b0,-10'd70,10'd70,-10'd70};
9'd235: value = {6'b0,-10'd70,10'd35,-10'd35};
9'd236: value = {6'b0,-10'd70,10'd0,10'd0};
9'd237: value = {6'b0,-10'd70,-10'd35,10'd35};
9'd238: value = {6'b0,-10'd70,-10'd70,10'd70};
9'd239: value = {6'b0,-10'd70,-10'd106,10'd106};
9'd240: value = {6'b0,-10'd106,10'd166,-10'd116};
9'd241: value = {6'b0,-10'd106,10'd131,-10'd81};
9'd242: value = {6'b0,-10'd106,10'd95,-10'd45};
9'd243: value = {6'b0,-10'd106,10'd60,-10'd10};
9'd244: value = {6'b0,-10'd106,10'd25,10'd25};
9'd245: value = {6'b0,-10'd106,-10'd10,10'd60};
9'd246: value = {6'b0,-10'd106,-10'd45,10'd95};
9'd247: value = {6'b0,-10'd106,-10'd81,10'd131};
9'd248: value = {6'b0,-10'd141,10'd191,-10'd91};
9'd249: value = {6'b0,-10'd141,10'd156,-10'd56};
9'd250: value = {6'b0,-10'd141,10'd120,-10'd20};
9'd251: value = {6'b0,-10'd141,10'd85,10'd14};
9'd252: value = {6'b0,-10'd141,10'd50,10'd50};
9'd253: value = {6'b0,-10'd141,10'd14,10'd85};
9'd254: value = {6'b0,-10'd141,-10'd20,10'd120};
9'd255: value = {6'b0,-10'd141,-10'd56,10'd156};
9'd256: value = {6'b0,10'd141,10'd41,-10'd241};
9'd257: value = {6'b0,10'd141,10'd6,-10'd206};
9'd258: value = {6'b0,10'd141,-10'd29,-10'd170};
9'd259: value = {6'b0,10'd141,-10'd64,-10'd135};
9'd260: value = {6'b0,10'd141,-10'd100,-10'd99};
9'd261: value = {6'b0,10'd141,-10'd135,-10'd64};
9'd262: value = {6'b0,10'd141,-10'd170,-10'd29};
9'd263: value = {6'b0,10'd141,-10'd206,10'd6};
9'd264: value = {6'b0,10'd106,10'd66,-10'd216};
9'd265: value = {6'b0,10'd106,10'd31,-10'd181};
9'd266: value = {6'b0,10'd106,-10'd4,-10'd145};
9'd267: value = {6'b0,10'd106,-10'd39,-10'd110};
9'd268: value = {6'b0,10'd106,-10'd75,-10'd74};
9'd269: value = {6'b0,10'd106,-10'd110,-10'd39};
9'd270: value = {6'b0,10'd106,-10'd145,-10'd4};
9'd271: value = {6'b0,10'd106,-10'd181,10'd31};
9'd272: value = {6'b0,10'd70,10'd91,-10'd191};
9'd273: value = {6'b0,10'd70,10'd56,-10'd156};
9'd274: value = {6'b0,10'd70,10'd20,-10'd120};
9'd275: value = {6'b0,10'd70,-10'd14,-10'd85};
9'd276: value = {6'b0,10'd70,-10'd50,-10'd49};
9'd277: value = {6'b0,10'd70,-10'd85,-10'd14};
9'd278: value = {6'b0,10'd70,-10'd120,10'd20};
9'd279: value = {6'b0,10'd70,-10'd156,10'd56};
9'd280: value = {6'b0,10'd35,10'd116,-10'd166};
9'd281: value = {6'b0,10'd35,10'd81,-10'd131};
9'd282: value = {6'b0,10'd35,10'd45,-10'd95};
9'd283: value = {6'b0,10'd35,10'd10,-10'd60};
9'd284: value = {6'b0,10'd35,-10'd25,-10'd24};
9'd285: value = {6'b0,10'd35,-10'd60,10'd10};
9'd286: value = {6'b0,10'd35,-10'd95,10'd45};
9'd287: value = {6'b0,10'd35,-10'd131,10'd81};
9'd288: value = {6'b0,10'd0,10'd141,-10'd141};
9'd289: value = {6'b0,10'd0,10'd106,-10'd106};
9'd290: value = {6'b0,10'd0,10'd70,-10'd70};
9'd291: value = {6'b0,10'd0,10'd35,-10'd35};
9'd292: value = {6'b0,10'd0,10'd0,10'd0};
9'd293: value = {6'b0,10'd0,-10'd35,10'd35};
9'd294: value = {6'b0,10'd0,-10'd70,10'd70};
9'd295: value = {6'b0,10'd0,-10'd106,10'd106};
9'd296: value = {6'b0,-10'd35,10'd166,-10'd116};
9'd297: value = {6'b0,-10'd35,10'd131,-10'd81};
9'd298: value = {6'b0,-10'd35,10'd95,-10'd45};
9'd299: value = {6'b0,-10'd35,10'd60,-10'd10};
9'd300: value = {6'b0,-10'd35,10'd25,10'd24};
9'd301: value = {6'b0,-10'd35,-10'd10,10'd60};
9'd302: value = {6'b0,-10'd35,-10'd45,10'd95};
9'd303: value = {6'b0,-10'd35,-10'd81,10'd131};
9'd304: value = {6'b0,-10'd70,10'd191,-10'd91};
9'd305: value = {6'b0,-10'd70,10'd156,-10'd56};
9'd306: value = {6'b0,-10'd70,10'd120,-10'd20};
9'd307: value = {6'b0,-10'd70,10'd85,10'd14};
9'd308: value = {6'b0,-10'd70,10'd50,10'd49};
9'd309: value = {6'b0,-10'd70,10'd14,10'd85};
9'd310: value = {6'b0,-10'd70,-10'd20,10'd120};
9'd311: value = {6'b0,-10'd70,-10'd56,10'd156};
9'd312: value = {6'b0,-10'd106,10'd216,-10'd66};
9'd313: value = {6'b0,-10'd106,10'd181,-10'd31};
9'd314: value = {6'b0,-10'd106,10'd145,10'd4};
9'd315: value = {6'b0,-10'd106,10'd110,10'd39};
9'd316: value = {6'b0,-10'd106,10'd75,10'd74};
9'd317: value = {6'b0,-10'd106,10'd39,10'd110};
9'd318: value = {6'b0,-10'd106,10'd4,10'd145};
9'd319: value = {6'b0,-10'd106,-10'd31,10'd181};
9'd320: value = {6'b0,10'd176,10'd66,-10'd216};
9'd321: value = {6'b0,10'd176,10'd31,-10'd181};
9'd322: value = {6'b0,10'd176,-10'd4,-10'd145};
9'd323: value = {6'b0,10'd176,-10'd39,-10'd110};
9'd324: value = {6'b0,10'd176,-10'd75,-10'd75};
9'd325: value = {6'b0,10'd176,-10'd110,-10'd39};
9'd326: value = {6'b0,10'd176,-10'd145,-10'd4};
9'd327: value = {6'b0,10'd176,-10'd181,10'd31};
9'd328: value = {6'b0,10'd141,10'd91,-10'd191};
9'd329: value = {6'b0,10'd141,10'd56,-10'd156};
9'd330: value = {6'b0,10'd141,10'd20,-10'd120};
9'd331: value = {6'b0,10'd141,-10'd14,-10'd85};
9'd332: value = {6'b0,10'd141,-10'd50,-10'd50};
9'd333: value = {6'b0,10'd141,-10'd85,-10'd14};
9'd334: value = {6'b0,10'd141,-10'd120,10'd20};
9'd335: value = {6'b0,10'd141,-10'd156,10'd56};
9'd336: value = {6'b0,10'd106,10'd116,-10'd166};
9'd337: value = {6'b0,10'd106,10'd81,-10'd131};
9'd338: value = {6'b0,10'd106,10'd45,-10'd95};
9'd339: value = {6'b0,10'd106,10'd10,-10'd60};
9'd340: value = {6'b0,10'd106,-10'd25,-10'd25};
9'd341: value = {6'b0,10'd106,-10'd60,10'd10};
9'd342: value = {6'b0,10'd106,-10'd95,10'd45};
9'd343: value = {6'b0,10'd106,-10'd131,10'd81};
9'd344: value = {6'b0,10'd70,10'd141,-10'd141};
9'd345: value = {6'b0,10'd70,10'd106,-10'd106};
9'd346: value = {6'b0,10'd70,10'd70,-10'd70};
9'd347: value = {6'b0,10'd70,10'd35,-10'd35};
9'd348: value = {6'b0,10'd70,-10'd0,-10'd0};
9'd349: value = {6'b0,10'd70,-10'd35,10'd35};
9'd350: value = {6'b0,10'd70,-10'd70,10'd70};
9'd351: value = {6'b0,10'd70,-10'd106,10'd106};
9'd352: value = {6'b0,10'd35,10'd166,-10'd116};
9'd353: value = {6'b0,10'd35,10'd131,-10'd81};
9'd354: value = {6'b0,10'd35,10'd95,-10'd45};
9'd355: value = {6'b0,10'd35,10'd60,-10'd10};
9'd356: value = {6'b0,10'd35,10'd24,10'd24};
9'd357: value = {6'b0,10'd35,-10'd10,10'd60};
9'd358: value = {6'b0,10'd35,-10'd45,10'd95};
9'd359: value = {6'b0,10'd35,-10'd81,10'd131};
9'd360: value = {6'b0,10'd0,10'd191,-10'd91};
9'd361: value = {6'b0,10'd0,10'd156,-10'd56};
9'd362: value = {6'b0,10'd0,10'd120,-10'd20};
9'd363: value = {6'b0,10'd0,10'd85,10'd14};
9'd364: value = {6'b0,10'd0,10'd50,10'd49};
9'd365: value = {6'b0,10'd0,10'd14,10'd85};
9'd366: value = {6'b0,10'd0,-10'd20,10'd120};
9'd367: value = {6'b0,10'd0,-10'd56,10'd156};
9'd368: value = {6'b0,-10'd35,10'd216,-10'd66};
9'd369: value = {6'b0,-10'd35,10'd181,-10'd31};
9'd370: value = {6'b0,-10'd35,10'd145,10'd4};
9'd371: value = {6'b0,-10'd35,10'd110,10'd39};
9'd372: value = {6'b0,-10'd35,10'd75,10'd74};
9'd373: value = {6'b0,-10'd35,10'd39,10'd110};
9'd374: value = {6'b0,-10'd35,10'd4,10'd145};
9'd375: value = {6'b0,-10'd35,-10'd31,10'd181};
9'd376: value = {6'b0,-10'd70,10'd241,-10'd41};
9'd377: value = {6'b0,-10'd70,10'd206,-10'd6};
9'd378: value = {6'b0,-10'd70,10'd170,10'd29};
9'd379: value = {6'b0,-10'd70,10'd135,10'd64};
9'd380: value = {6'b0,-10'd70,10'd100,10'd99};
9'd381: value = {6'b0,-10'd70,10'd64,10'd135};
9'd382: value = {6'b0,-10'd70,10'd29,10'd170};
9'd383: value = {6'b0,-10'd70,-10'd6,10'd206};
9'd384: value = {6'b0,10'd212,10'd91,-10'd191};
9'd385: value = {6'b0,10'd212,10'd56,-10'd156};
9'd386: value = {6'b0,10'd212,10'd20,-10'd120};
9'd387: value = {6'b0,10'd212,-10'd14,-10'd85};
9'd388: value = {6'b0,10'd212,-10'd50,-10'd50};
9'd389: value = {6'b0,10'd212,-10'd85,-10'd14};
9'd390: value = {6'b0,10'd212,-10'd120,10'd20};
9'd391: value = {6'b0,10'd212,-10'd156,10'd56};
9'd392: value = {6'b0,10'd176,10'd116,-10'd166};
9'd393: value = {6'b0,10'd176,10'd81,-10'd131};
9'd394: value = {6'b0,10'd176,10'd45,-10'd95};
9'd395: value = {6'b0,10'd176,10'd10,-10'd60};
9'd396: value = {6'b0,10'd176,-10'd25,-10'd25};
9'd397: value = {6'b0,10'd176,-10'd60,10'd10};
9'd398: value = {6'b0,10'd176,-10'd95,10'd45};
9'd399: value = {6'b0,10'd176,-10'd131,10'd81};
9'd400: value = {6'b0,10'd141,10'd141,-10'd141};
9'd401: value = {6'b0,10'd141,10'd106,-10'd106};
9'd402: value = {6'b0,10'd141,10'd70,-10'd70};
9'd403: value = {6'b0,10'd141,10'd35,-10'd35};
9'd404: value = {6'b0,10'd141,-10'd0,-10'd0};
9'd405: value = {6'b0,10'd141,-10'd35,10'd35};
9'd406: value = {6'b0,10'd141,-10'd70,10'd70};
9'd407: value = {6'b0,10'd141,-10'd106,10'd106};
9'd408: value = {6'b0,10'd106,10'd166,-10'd116};
9'd409: value = {6'b0,10'd106,10'd131,-10'd81};
9'd410: value = {6'b0,10'd106,10'd95,-10'd45};
9'd411: value = {6'b0,10'd106,10'd60,-10'd10};
9'd412: value = {6'b0,10'd106,10'd24,10'd24};
9'd413: value = {6'b0,10'd106,-10'd10,10'd60};
9'd414: value = {6'b0,10'd106,-10'd45,10'd95};
9'd415: value = {6'b0,10'd106,-10'd81,10'd131};
9'd416: value = {6'b0,10'd70,10'd191,-10'd91};
9'd417: value = {6'b0,10'd70,10'd156,-10'd56};
9'd418: value = {6'b0,10'd70,10'd120,-10'd20};
9'd419: value = {6'b0,10'd70,10'd85,10'd14};
9'd420: value = {6'b0,10'd70,10'd49,10'd49};
9'd421: value = {6'b0,10'd70,10'd14,10'd85};
9'd422: value = {6'b0,10'd70,-10'd20,10'd120};
9'd423: value = {6'b0,10'd70,-10'd56,10'd156};
9'd424: value = {6'b0,10'd35,10'd216,-10'd66};
9'd425: value = {6'b0,10'd35,10'd181,-10'd31};
9'd426: value = {6'b0,10'd35,10'd145,10'd4};
9'd427: value = {6'b0,10'd35,10'd110,10'd39};
9'd428: value = {6'b0,10'd35,10'd75,10'd74};
9'd429: value = {6'b0,10'd35,10'd39,10'd110};
9'd430: value = {6'b0,10'd35,10'd4,10'd145};
9'd431: value = {6'b0,10'd35,-10'd31,10'd181};
9'd432: value = {6'b0,10'd0,10'd241,-10'd41};
9'd433: value = {6'b0,10'd0,10'd206,-10'd6};
9'd434: value = {6'b0,10'd0,10'd170,10'd29};
9'd435: value = {6'b0,10'd0,10'd135,10'd64};
9'd436: value = {6'b0,10'd0,10'd100,10'd99};
9'd437: value = {6'b0,10'd0,10'd64,10'd135};
9'd438: value = {6'b0,10'd0,10'd29,10'd170};
9'd439: value = {6'b0,10'd0,-10'd6,10'd206};
9'd440: value = {6'b0,-10'd35,10'd266,-10'd16};
9'd441: value = {6'b0,-10'd35,10'd231,10'd18};
9'd442: value = {6'b0,-10'd35,10'd195,10'd54};
9'd443: value = {6'b0,-10'd35,10'd160,10'd89};
9'd444: value = {6'b0,-10'd35,10'd125,10'd124};
9'd445: value = {6'b0,-10'd35,10'd89,10'd160};
9'd446: value = {6'b0,-10'd35,10'd54,10'd195};
9'd447: value = {6'b0,-10'd35,10'd18,10'd231};
9'd448: value = {6'b0,10'd247,10'd116,-10'd166};
9'd449: value = {6'b0,10'd247,10'd81,-10'd131};
9'd450: value = {6'b0,10'd247,10'd45,-10'd95};
9'd451: value = {6'b0,10'd247,10'd10,-10'd60};
9'd452: value = {6'b0,10'd247,-10'd25,-10'd25};
9'd453: value = {6'b0,10'd247,-10'd60,10'd10};
9'd454: value = {6'b0,10'd247,-10'd95,10'd45};
9'd455: value = {6'b0,10'd247,-10'd131,10'd81};
9'd456: value = {6'b0,10'd212,10'd141,-10'd141};
9'd457: value = {6'b0,10'd212,10'd106,-10'd106};
9'd458: value = {6'b0,10'd212,10'd70,-10'd70};
9'd459: value = {6'b0,10'd212,10'd35,-10'd35};
9'd460: value = {6'b0,10'd212,-10'd0,-10'd0};
9'd461: value = {6'b0,10'd212,-10'd35,10'd35};
9'd462: value = {6'b0,10'd212,-10'd70,10'd70};
9'd463: value = {6'b0,10'd212,-10'd106,10'd106};
9'd464: value = {6'b0,10'd176,10'd166,-10'd116};
9'd465: value = {6'b0,10'd176,10'd131,-10'd81};
9'd466: value = {6'b0,10'd176,10'd95,-10'd45};
9'd467: value = {6'b0,10'd176,10'd60,-10'd10};
9'd468: value = {6'b0,10'd176,10'd24,10'd24};
9'd469: value = {6'b0,10'd176,-10'd10,10'd60};
9'd470: value = {6'b0,10'd176,-10'd45,10'd95};
9'd471: value = {6'b0,10'd176,-10'd81,10'd131};
9'd472: value = {6'b0,10'd141,10'd191,-10'd91};
9'd473: value = {6'b0,10'd141,10'd156,-10'd56};
9'd474: value = {6'b0,10'd141,10'd120,-10'd20};
9'd475: value = {6'b0,10'd141,10'd85,10'd14};
9'd476: value = {6'b0,10'd141,10'd49,10'd49};
9'd477: value = {6'b0,10'd141,10'd14,10'd85};
9'd478: value = {6'b0,10'd141,-10'd20,10'd120};
9'd479: value = {6'b0,10'd141,-10'd56,10'd156};
9'd480: value = {6'b0,10'd106,10'd216,-10'd66};
9'd481: value = {6'b0,10'd106,10'd181,-10'd31};
9'd482: value = {6'b0,10'd106,10'd145,10'd4};
9'd483: value = {6'b0,10'd106,10'd110,10'd39};
9'd484: value = {6'b0,10'd106,10'd74,10'd74};
9'd485: value = {6'b0,10'd106,10'd39,10'd110};
9'd486: value = {6'b0,10'd106,10'd4,10'd145};
9'd487: value = {6'b0,10'd106,-10'd31,10'd181};
9'd488: value = {6'b0,10'd70,10'd241,-10'd41};
9'd489: value = {6'b0,10'd70,10'd206,-10'd6};
9'd490: value = {6'b0,10'd70,10'd170,10'd29};
9'd491: value = {6'b0,10'd70,10'd135,10'd64};
9'd492: value = {6'b0,10'd70,10'd100,10'd99};
9'd493: value = {6'b0,10'd70,10'd64,10'd135};
9'd494: value = {6'b0,10'd70,10'd29,10'd170};
9'd495: value = {6'b0,10'd70,-10'd6,10'd206};
9'd496: value = {6'b0,10'd35,10'd266,-10'd16};
9'd497: value = {6'b0,10'd35,10'd231,10'd18};
9'd498: value = {6'b0,10'd35,10'd195,10'd54};
9'd499: value = {6'b0,10'd35,10'd160,10'd89};
9'd500: value = {6'b0,10'd35,10'd125,10'd124};
9'd501: value = {6'b0,10'd35,10'd89,10'd160};
9'd502: value = {6'b0,10'd35,10'd54,10'd195};
9'd503: value = {6'b0,10'd35,10'd18,10'd231};
9'd504: value = {6'b0,10'd0,10'd291,10'd8};
9'd505: value = {6'b0,10'd0,10'd256,10'd43};
9'd506: value = {6'b0,10'd0,10'd220,10'd79};
9'd507: value = {6'b0,10'd0,10'd185,10'd114};
9'd508: value = {6'b0,10'd0,10'd150,10'd149};
9'd509: value = {6'b0,10'd0,10'd114,10'd185};
9'd510: value = {6'b0,10'd0,10'd79,10'd220};
9'd511: value = {6'b0,10'd0,10'd43,10'd256};
			default: value = 0;
		endcase
endmodule
